-- nios_ii_base.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_ii_base is
	port (
		clk_clk            : in    std_logic                     := '0';             --         clk.clk
		hex_3_HEX0         : out   std_logic_vector(6 downto 0);                     --       hex_3.HEX0
		hex_3_HEX1         : out   std_logic_vector(6 downto 0);                     --            .HEX1
		hex_3_HEX2         : out   std_logic_vector(6 downto 0);                     --            .HEX2
		hex_3_HEX3         : out   std_logic_vector(6 downto 0);                     --            .HEX3
		hex_7_HEX4         : out   std_logic_vector(6 downto 0);                     --       hex_7.HEX4
		hex_7_HEX5         : out   std_logic_vector(6 downto 0);                     --            .HEX5
		hex_7_HEX6         : out   std_logic_vector(6 downto 0);                     --            .HEX6
		hex_7_HEX7         : out   std_logic_vector(6 downto 0);                     --            .HEX7
		lcd_DATA           : inout std_logic_vector(7 downto 0)  := (others => '0'); --         lcd.DATA
		lcd_ON             : out   std_logic;                                        --            .ON
		lcd_BLON           : out   std_logic;                                        --            .BLON
		lcd_EN             : out   std_logic;                                        --            .EN
		lcd_RS             : out   std_logic;                                        --            .RS
		lcd_RW             : out   std_logic;                                        --            .RW
		leds_green_export  : out   std_logic_vector(8 downto 0);                     --  leds_green.export
		leds_red_export    : out   std_logic_vector(17 downto 0);                    --    leds_red.export
		pushbuttons_export : in    std_logic_vector(3 downto 0)  := (others => '0'); -- pushbuttons.export
		reset_reset_n      : in    std_logic                     := '0';             --       reset.reset_n
		sw_sliders_export  : in    std_logic_vector(17 downto 0) := (others => '0'); --  sw_sliders.export
		vga_CLK            : out   std_logic;                                        --         vga.CLK
		vga_HS             : out   std_logic;                                        --            .HS
		vga_VS             : out   std_logic;                                        --            .VS
		vga_BLANK          : out   std_logic;                                        --            .BLANK
		vga_SYNC           : out   std_logic;                                        --            .SYNC
		vga_R              : out   std_logic_vector(7 downto 0);                     --            .R
		vga_G              : out   std_logic_vector(7 downto 0);                     --            .G
		vga_B              : out   std_logic_vector(7 downto 0)                      --            .B
	);
end entity nios_ii_base;

architecture rtl of nios_ii_base is
	component nios_ii_base_HEX_3 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			HEX0       : out std_logic_vector(6 downto 0);                     -- export
			HEX1       : out std_logic_vector(6 downto 0);                     -- export
			HEX2       : out std_logic_vector(6 downto 0);                     -- export
			HEX3       : out std_logic_vector(6 downto 0)                      -- export
		);
	end component nios_ii_base_HEX_3;

	component nios_ii_base_HEX_7 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			HEX4       : out std_logic_vector(6 downto 0);                     -- export
			HEX5       : out std_logic_vector(6 downto 0);                     -- export
			HEX6       : out std_logic_vector(6 downto 0);                     -- export
			HEX7       : out std_logic_vector(6 downto 0)                      -- export
		);
	end component nios_ii_base_HEX_7;

	component nios_ii_base_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_ii_base_JTAG_UART;

	component nios_ii_base_LCD is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component nios_ii_base_LCD;

	component nios_ii_base_LEDS_GREEN is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDG       : out std_logic_vector(8 downto 0)                      -- export
		);
	end component nios_ii_base_LEDS_GREEN;

	component nios_ii_base_LEDS_RED is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDR       : out std_logic_vector(17 downto 0)                     -- export
		);
	end component nios_ii_base_LEDS_RED;

	component nios_ii_base_NIOS_II_Processor is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_ii_base_NIOS_II_Processor;

	component nios_ii_base_OnChip_Memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(63 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_ii_base_OnChip_Memory;

	component nios_ii_base_Pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			KEY        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_ii_base_Pushbuttons;

	component nios_ii_base_SW_SLIDERS is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			SW         : in  std_logic_vector(17 downto 0) := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_ii_base_SW_SLIDERS;

	component nios_ii_base_VGA_Char_Buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component nios_ii_base_VGA_Char_Buffer;

	component nios_ii_base_VGA_Controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_ii_base_VGA_Controller;

	component nios_ii_base_VGA_Dual_Clock_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component nios_ii_base_VGA_Dual_Clock_FIFO;

	component nios_ii_base_VGA_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component nios_ii_base_VGA_PLL;

	component nios_ii_base_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_ii_base_timer_0;

	component nios_ii_base_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			NIOS_II_Processor_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			VGA_Char_Buffer_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			NIOS_II_Processor_data_master_address                : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NIOS_II_Processor_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			NIOS_II_Processor_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS_II_Processor_data_master_read                   : in  std_logic                     := 'X';             -- read
			NIOS_II_Processor_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_II_Processor_data_master_write                  : in  std_logic                     := 'X';             -- write
			NIOS_II_Processor_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS_II_Processor_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			NIOS_II_Processor_instruction_master_address         : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NIOS_II_Processor_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			NIOS_II_Processor_instruction_master_read            : in  std_logic                     := 'X';             -- read
			NIOS_II_Processor_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			HEX_3_avalon_parallel_port_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			HEX_3_avalon_parallel_port_slave_write               : out std_logic;                                        -- write
			HEX_3_avalon_parallel_port_slave_read                : out std_logic;                                        -- read
			HEX_3_avalon_parallel_port_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_3_avalon_parallel_port_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_3_avalon_parallel_port_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			HEX_3_avalon_parallel_port_slave_chipselect          : out std_logic;                                        -- chipselect
			HEX_7_avalon_parallel_port_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			HEX_7_avalon_parallel_port_slave_write               : out std_logic;                                        -- write
			HEX_7_avalon_parallel_port_slave_read                : out std_logic;                                        -- read
			HEX_7_avalon_parallel_port_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX_7_avalon_parallel_port_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			HEX_7_avalon_parallel_port_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			HEX_7_avalon_parallel_port_slave_chipselect          : out std_logic;                                        -- chipselect
			JTAG_UART_avalon_jtag_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                    : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                     : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect               : out std_logic;                                        -- chipselect
			LCD_avalon_lcd_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			LCD_avalon_lcd_slave_write                           : out std_logic;                                        -- write
			LCD_avalon_lcd_slave_read                            : out std_logic;                                        -- read
			LCD_avalon_lcd_slave_readdata                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			LCD_avalon_lcd_slave_writedata                       : out std_logic_vector(7 downto 0);                     -- writedata
			LCD_avalon_lcd_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			LCD_avalon_lcd_slave_chipselect                      : out std_logic;                                        -- chipselect
			LEDS_GREEN_avalon_parallel_port_slave_address        : out std_logic_vector(1 downto 0);                     -- address
			LEDS_GREEN_avalon_parallel_port_slave_write          : out std_logic;                                        -- write
			LEDS_GREEN_avalon_parallel_port_slave_read           : out std_logic;                                        -- read
			LEDS_GREEN_avalon_parallel_port_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDS_GREEN_avalon_parallel_port_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			LEDS_GREEN_avalon_parallel_port_slave_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			LEDS_GREEN_avalon_parallel_port_slave_chipselect     : out std_logic;                                        -- chipselect
			LEDS_RED_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			LEDS_RED_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			LEDS_RED_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			LEDS_RED_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDS_RED_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			LEDS_RED_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			LEDS_RED_avalon_parallel_port_slave_chipselect       : out std_logic;                                        -- chipselect
			NIOS_II_Processor_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			NIOS_II_Processor_debug_mem_slave_write              : out std_logic;                                        -- write
			NIOS_II_Processor_debug_mem_slave_read               : out std_logic;                                        -- read
			NIOS_II_Processor_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS_II_Processor_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS_II_Processor_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS_II_Processor_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			NIOS_II_Processor_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			OnChip_Memory_s1_address                             : out std_logic_vector(14 downto 0);                    -- address
			OnChip_Memory_s1_write                               : out std_logic;                                        -- write
			OnChip_Memory_s1_readdata                            : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			OnChip_Memory_s1_writedata                           : out std_logic_vector(63 downto 0);                    -- writedata
			OnChip_Memory_s1_byteenable                          : out std_logic_vector(7 downto 0);                     -- byteenable
			OnChip_Memory_s1_chipselect                          : out std_logic;                                        -- chipselect
			OnChip_Memory_s1_clken                               : out std_logic;                                        -- clken
			Pushbuttons_avalon_parallel_port_slave_address       : out std_logic_vector(1 downto 0);                     -- address
			Pushbuttons_avalon_parallel_port_slave_write         : out std_logic;                                        -- write
			Pushbuttons_avalon_parallel_port_slave_read          : out std_logic;                                        -- read
			Pushbuttons_avalon_parallel_port_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pushbuttons_avalon_parallel_port_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			Pushbuttons_avalon_parallel_port_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			Pushbuttons_avalon_parallel_port_slave_chipselect    : out std_logic;                                        -- chipselect
			SW_SLIDERS_avalon_parallel_port_slave_address        : out std_logic_vector(1 downto 0);                     -- address
			SW_SLIDERS_avalon_parallel_port_slave_write          : out std_logic;                                        -- write
			SW_SLIDERS_avalon_parallel_port_slave_read           : out std_logic;                                        -- read
			SW_SLIDERS_avalon_parallel_port_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SW_SLIDERS_avalon_parallel_port_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			SW_SLIDERS_avalon_parallel_port_slave_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			SW_SLIDERS_avalon_parallel_port_slave_chipselect     : out std_logic;                                        -- chipselect
			timer_0_s1_address                                   : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                     : out std_logic;                                        -- write
			timer_0_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                : out std_logic;                                        -- chipselect
			timer_1_s1_address                                   : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                     : out std_logic;                                        -- write
			timer_1_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                                : out std_logic;                                        -- chipselect
			VGA_Char_Buffer_avalon_char_buffer_slave_address     : out std_logic_vector(12 downto 0);                    -- address
			VGA_Char_Buffer_avalon_char_buffer_slave_write       : out std_logic;                                        -- write
			VGA_Char_Buffer_avalon_char_buffer_slave_read        : out std_logic;                                        -- read
			VGA_Char_Buffer_avalon_char_buffer_slave_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			VGA_Char_Buffer_avalon_char_buffer_slave_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			VGA_Char_Buffer_avalon_char_buffer_slave_byteenable  : out std_logic_vector(0 downto 0);                     -- byteenable
			VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			VGA_Char_Buffer_avalon_char_buffer_slave_chipselect  : out std_logic;                                        -- chipselect
			VGA_Char_Buffer_avalon_char_control_slave_address    : out std_logic_vector(0 downto 0);                     -- address
			VGA_Char_Buffer_avalon_char_control_slave_write      : out std_logic;                                        -- write
			VGA_Char_Buffer_avalon_char_control_slave_read       : out std_logic;                                        -- read
			VGA_Char_Buffer_avalon_char_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VGA_Char_Buffer_avalon_char_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_Char_Buffer_avalon_char_control_slave_byteenable : out std_logic_vector(3 downto 0);                     -- byteenable
			VGA_Char_Buffer_avalon_char_control_slave_chipselect : out std_logic                                         -- chipselect
		);
	end component nios_ii_base_mm_interconnect_0;

	component nios_ii_base_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_ii_base_irq_mapper;

	component nios_ii_base_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_ii_base_rst_controller;

	component nios_ii_base_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_ii_base_rst_controller_001;

	signal vga_char_buffer_avalon_char_source_valid                               : std_logic;                     -- VGA_Char_Buffer:stream_valid -> VGA_Dual_Clock_FIFO:stream_in_valid
	signal vga_char_buffer_avalon_char_source_data                                : std_logic_vector(29 downto 0); -- VGA_Char_Buffer:stream_data -> VGA_Dual_Clock_FIFO:stream_in_data
	signal vga_char_buffer_avalon_char_source_ready                               : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_in_ready -> VGA_Char_Buffer:stream_ready
	signal vga_char_buffer_avalon_char_source_startofpacket                       : std_logic;                     -- VGA_Char_Buffer:stream_startofpacket -> VGA_Dual_Clock_FIFO:stream_in_startofpacket
	signal vga_char_buffer_avalon_char_source_endofpacket                         : std_logic;                     -- VGA_Char_Buffer:stream_endofpacket -> VGA_Dual_Clock_FIFO:stream_in_endofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_valid                      : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_data                       : std_logic_vector(29 downto 0); -- VGA_Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_ready                      : std_logic;                     -- VGA_Controller:ready -> VGA_Dual_Clock_FIFO:stream_out_ready
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket              : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket                : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	signal vga_pll_vga_clk_clk                                                    : std_logic;                     -- VGA_PLL:vga_clk_clk -> [VGA_Controller:clk, VGA_Dual_Clock_FIFO:clk_stream_out, rst_controller_002:clk]
	signal nios_ii_processor_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_data_master_readdata -> NIOS_II_Processor:d_readdata
	signal nios_ii_processor_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_data_master_waitrequest -> NIOS_II_Processor:d_waitrequest
	signal nios_ii_processor_data_master_debugaccess                              : std_logic;                     -- NIOS_II_Processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_II_Processor_data_master_debugaccess
	signal nios_ii_processor_data_master_address                                  : std_logic_vector(19 downto 0); -- NIOS_II_Processor:d_address -> mm_interconnect_0:NIOS_II_Processor_data_master_address
	signal nios_ii_processor_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- NIOS_II_Processor:d_byteenable -> mm_interconnect_0:NIOS_II_Processor_data_master_byteenable
	signal nios_ii_processor_data_master_read                                     : std_logic;                     -- NIOS_II_Processor:d_read -> mm_interconnect_0:NIOS_II_Processor_data_master_read
	signal nios_ii_processor_data_master_write                                    : std_logic;                     -- NIOS_II_Processor:d_write -> mm_interconnect_0:NIOS_II_Processor_data_master_write
	signal nios_ii_processor_data_master_writedata                                : std_logic_vector(31 downto 0); -- NIOS_II_Processor:d_writedata -> mm_interconnect_0:NIOS_II_Processor_data_master_writedata
	signal nios_ii_processor_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_instruction_master_readdata -> NIOS_II_Processor:i_readdata
	signal nios_ii_processor_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_instruction_master_waitrequest -> NIOS_II_Processor:i_waitrequest
	signal nios_ii_processor_instruction_master_address                           : std_logic_vector(19 downto 0); -- NIOS_II_Processor:i_address -> mm_interconnect_0:NIOS_II_Processor_instruction_master_address
	signal nios_ii_processor_instruction_master_read                              : std_logic;                     -- NIOS_II_Processor:i_read -> mm_interconnect_0:NIOS_II_Processor_instruction_master_read
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_chipselect  : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_chipselect -> VGA_Char_Buffer:buf_chipselect
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_readdata    : std_logic_vector(7 downto 0);  -- VGA_Char_Buffer:buf_readdata -> mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_readdata
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_waitrequest : std_logic;                     -- VGA_Char_Buffer:buf_waitrequest -> mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_address     : std_logic_vector(12 downto 0); -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_address -> VGA_Char_Buffer:buf_address
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_read        : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_read -> VGA_Char_Buffer:buf_read
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_byteenable  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_byteenable -> VGA_Char_Buffer:buf_byteenable
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_write       : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_write -> VGA_Char_Buffer:buf_write
	signal mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_buffer_slave_writedata -> VGA_Char_Buffer:buf_writedata
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_chipselect : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_chipselect -> VGA_Char_Buffer:ctrl_chipselect
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_readdata   : std_logic_vector(31 downto 0); -- VGA_Char_Buffer:ctrl_readdata -> mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_readdata
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_address    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_address -> VGA_Char_Buffer:ctrl_address
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_read       : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_read -> VGA_Char_Buffer:ctrl_read
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_byteenable -> VGA_Char_Buffer:ctrl_byteenable
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_write      : std_logic;                     -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_write -> VGA_Char_Buffer:ctrl_write
	signal mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_Char_Buffer_avalon_char_control_slave_writedata -> VGA_Char_Buffer:ctrl_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect               : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                 : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest              : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                     : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                    : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_lcd_avalon_lcd_slave_chipselect                      : std_logic;                     -- mm_interconnect_0:LCD_avalon_lcd_slave_chipselect -> LCD:chipselect
	signal mm_interconnect_0_lcd_avalon_lcd_slave_readdata                        : std_logic_vector(7 downto 0);  -- LCD:readdata -> mm_interconnect_0:LCD_avalon_lcd_slave_readdata
	signal mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest                     : std_logic;                     -- LCD:waitrequest -> mm_interconnect_0:LCD_avalon_lcd_slave_waitrequest
	signal mm_interconnect_0_lcd_avalon_lcd_slave_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:LCD_avalon_lcd_slave_address -> LCD:address
	signal mm_interconnect_0_lcd_avalon_lcd_slave_read                            : std_logic;                     -- mm_interconnect_0:LCD_avalon_lcd_slave_read -> LCD:read
	signal mm_interconnect_0_lcd_avalon_lcd_slave_write                           : std_logic;                     -- mm_interconnect_0:LCD_avalon_lcd_slave_write -> LCD:write
	signal mm_interconnect_0_lcd_avalon_lcd_slave_writedata                       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:LCD_avalon_lcd_slave_writedata -> LCD:writedata
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_chipselect     : std_logic;                     -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_chipselect -> SW_SLIDERS:chipselect
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_readdata       : std_logic_vector(31 downto 0); -- SW_SLIDERS:readdata -> mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_address -> SW_SLIDERS:address
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_read           : std_logic;                     -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_read -> SW_SLIDERS:read
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_byteenable -> SW_SLIDERS:byteenable
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_write          : std_logic;                     -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_write -> SW_SLIDERS:write
	signal mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:SW_SLIDERS_avalon_parallel_port_slave_writedata -> SW_SLIDERS:writedata
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_chipselect     : std_logic;                     -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_chipselect -> LEDS_GREEN:chipselect
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_readdata       : std_logic_vector(31 downto 0); -- LEDS_GREEN:readdata -> mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_address -> LEDS_GREEN:address
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_read           : std_logic;                     -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_read -> LEDS_GREEN:read
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_byteenable -> LEDS_GREEN:byteenable
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_write          : std_logic;                     -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_write -> LEDS_GREEN:write
	signal mm_interconnect_0_leds_green_avalon_parallel_port_slave_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDS_GREEN_avalon_parallel_port_slave_writedata -> LEDS_GREEN:writedata
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_chipselect       : std_logic;                     -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_chipselect -> LEDS_RED:chipselect
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_readdata         : std_logic_vector(31 downto 0); -- LEDS_RED:readdata -> mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_address          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_address -> LEDS_RED:address
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_read             : std_logic;                     -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_read -> LEDS_RED:read
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_byteenable -> LEDS_RED:byteenable
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_write            : std_logic;                     -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_write -> LEDS_RED:write
	signal mm_interconnect_0_leds_red_avalon_parallel_port_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDS_RED_avalon_parallel_port_slave_writedata -> LEDS_RED:writedata
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_chipselect          : std_logic;                     -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_chipselect -> HEX_3:chipselect
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_readdata            : std_logic_vector(31 downto 0); -- HEX_3:readdata -> mm_interconnect_0:HEX_3_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_address -> HEX_3:address
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_read                : std_logic;                     -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_read -> HEX_3:read
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_byteenable -> HEX_3:byteenable
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_write               : std_logic;                     -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_write -> HEX_3:write
	signal mm_interconnect_0_hex_3_avalon_parallel_port_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_3_avalon_parallel_port_slave_writedata -> HEX_3:writedata
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_chipselect          : std_logic;                     -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_chipselect -> HEX_7:chipselect
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_readdata            : std_logic_vector(31 downto 0); -- HEX_7:readdata -> mm_interconnect_0:HEX_7_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_address -> HEX_7:address
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_read                : std_logic;                     -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_read -> HEX_7:read
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_byteenable -> HEX_7:byteenable
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_write               : std_logic;                     -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_write -> HEX_7:write
	signal mm_interconnect_0_hex_7_avalon_parallel_port_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX_7_avalon_parallel_port_slave_writedata -> HEX_7:writedata
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect    : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_chipselect -> Pushbuttons:chipselect
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata      : std_logic_vector(31 downto 0); -- Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_address -> Pushbuttons:address
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read          : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_read -> Pushbuttons:read
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_byteenable -> Pushbuttons:byteenable
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write         : std_logic;                     -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_write -> Pushbuttons:write
	signal mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_writedata -> Pushbuttons:writedata
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- NIOS_II_Processor:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest        : std_logic;                     -- NIOS_II_Processor:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_debugaccess -> NIOS_II_Processor:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_address -> NIOS_II_Processor:debug_mem_slave_address
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_read -> NIOS_II_Processor:debug_mem_slave_read
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_byteenable -> NIOS_II_Processor:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_write -> NIOS_II_Processor:debug_mem_slave_write
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_writedata -> NIOS_II_Processor:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_chipselect -> OnChip_Memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                            : std_logic_vector(63 downto 0); -- OnChip_Memory:readdata -> mm_interconnect_0:OnChip_Memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                             : std_logic_vector(14 downto 0); -- mm_interconnect_0:OnChip_Memory_s1_address -> OnChip_Memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:OnChip_Memory_s1_byteenable -> OnChip_Memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                               : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_write -> OnChip_Memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                           : std_logic_vector(63 downto 0); -- mm_interconnect_0:OnChip_Memory_s1_writedata -> OnChip_Memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                               : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_clken -> OnChip_Memory:clken
	signal mm_interconnect_0_timer_0_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                  : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                     : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                                  : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                                     : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal irq_mapper_receiver0_irq                                               : std_logic;                     -- SW_SLIDERS:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                               : std_logic;                     -- Pushbuttons:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                               : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                               : std_logic;                     -- timer_0:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                               : std_logic;                     -- timer_1:irq -> irq_mapper:receiver4_irq
	signal nios_ii_processor_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS_II_Processor:irq
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [HEX_3:reset, HEX_7:reset, LCD:reset, LEDS_GREEN:reset, LEDS_RED:reset, OnChip_Memory:reset, Pushbuttons:reset, SW_SLIDERS:reset, irq_mapper:reset, mm_interconnect_0:NIOS_II_Processor_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                     : std_logic;                     -- rst_controller:reset_req -> [NIOS_II_Processor:reset_req, OnChip_Memory:reset_req, rst_translator:reset_req_in]
	signal nios_ii_processor_debug_reset_request_reset                            : std_logic;                     -- NIOS_II_Processor:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                                     : std_logic;                     -- rst_controller_001:reset_out -> [VGA_Char_Buffer:reset, VGA_Dual_Clock_FIFO:reset_stream_in, VGA_PLL:ref_reset_reset, mm_interconnect_0:VGA_Char_Buffer_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                                     : std_logic;                     -- rst_controller_002:reset_out -> [VGA_Controller:reset, VGA_Dual_Clock_FIFO:reset_stream_out]
	signal vga_pll_reset_source_reset                                             : std_logic;                     -- VGA_PLL:reset_source_reset -> rst_controller_002:reset_in0
	signal reset_reset_n_ports_inv                                                : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_UART:rst_n, NIOS_II_Processor:reset_n, timer_0:reset_n, timer_1:reset_n]

begin

	hex_3 : component nios_ii_base_HEX_3
		port map (
			clk        => clk_clk,                                                       --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                --                      reset.reset
			address    => mm_interconnect_0_hex_3_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_hex_3_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_hex_3_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_hex_3_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_hex_3_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_hex_3_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_hex_3_avalon_parallel_port_slave_readdata,   --                           .readdata
			HEX0       => hex_3_HEX0,                                                    --         external_interface.export
			HEX1       => hex_3_HEX1,                                                    --                           .export
			HEX2       => hex_3_HEX2,                                                    --                           .export
			HEX3       => hex_3_HEX3                                                     --                           .export
		);

	hex_7 : component nios_ii_base_HEX_7
		port map (
			clk        => clk_clk,                                                       --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                --                      reset.reset
			address    => mm_interconnect_0_hex_7_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_hex_7_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_hex_7_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_hex_7_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_hex_7_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_hex_7_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_hex_7_avalon_parallel_port_slave_readdata,   --                           .readdata
			HEX4       => hex_7_HEX4,                                                    --         external_interface.export
			HEX5       => hex_7_HEX5,                                                    --                           .export
			HEX6       => hex_7_HEX6,                                                    --                           .export
			HEX7       => hex_7_HEX7                                                     --                           .export
		);

	jtag_uart : component nios_ii_base_JTAG_UART
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                       --               irq.irq
		);

	lcd : component nios_ii_base_LCD
		port map (
			clk         => clk_clk,                                            --                clk.clk
			reset       => rst_controller_reset_out_reset,                     --              reset.reset
			address     => mm_interconnect_0_lcd_avalon_lcd_slave_address(0),  --   avalon_lcd_slave.address
			chipselect  => mm_interconnect_0_lcd_avalon_lcd_slave_chipselect,  --                   .chipselect
			read        => mm_interconnect_0_lcd_avalon_lcd_slave_read,        --                   .read
			write       => mm_interconnect_0_lcd_avalon_lcd_slave_write,       --                   .write
			writedata   => mm_interconnect_0_lcd_avalon_lcd_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_lcd_avalon_lcd_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest, --                   .waitrequest
			LCD_DATA    => lcd_DATA,                                           -- external_interface.export
			LCD_ON      => lcd_ON,                                             --                   .export
			LCD_BLON    => lcd_BLON,                                           --                   .export
			LCD_EN      => lcd_EN,                                             --                   .export
			LCD_RS      => lcd_RS,                                             --                   .export
			LCD_RW      => lcd_RW                                              --                   .export
		);

	leds_green : component nios_ii_base_LEDS_GREEN
		port map (
			clk        => clk_clk,                                                            --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                     --                      reset.reset
			address    => mm_interconnect_0_leds_green_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_leds_green_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_leds_green_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_leds_green_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_leds_green_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_leds_green_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_leds_green_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDG       => leds_green_export                                                   --         external_interface.export
		);

	leds_red : component nios_ii_base_LEDS_RED
		port map (
			clk        => clk_clk,                                                          --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                   --                      reset.reset
			address    => mm_interconnect_0_leds_red_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_leds_red_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_leds_red_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_leds_red_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_leds_red_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_leds_red_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_leds_red_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDR       => leds_red_export                                                   --         external_interface.export
		);

	nios_ii_processor : component nios_ii_base_NIOS_II_Processor
		port map (
			clk                                 => clk_clk,                                                         --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                        --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                              --                          .reset_req
			d_address                           => nios_ii_processor_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_ii_processor_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_ii_processor_data_master_read,                              --                          .read
			d_readdata                          => nios_ii_processor_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_ii_processor_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_ii_processor_data_master_write,                             --                          .write
			d_writedata                         => nios_ii_processor_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_ii_processor_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_ii_processor_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_ii_processor_instruction_master_read,                       --                          .read
			i_readdata                          => nios_ii_processor_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_ii_processor_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_ii_processor_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_ii_processor_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_ii_processor_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_ii_processor_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_ii_processor_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                             -- custom_instruction_master.readra
		);

	onchip_memory : component nios_ii_base_OnChip_Memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	pushbuttons : component nios_ii_base_Pushbuttons
		port map (
			clk        => clk_clk,                                                             --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                      --                      reset.reset
			address    => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata,   --                           .readdata
			KEY        => pushbuttons_export,                                                  --         external_interface.export
			irq        => irq_mapper_receiver1_irq                                             --                  interrupt.irq
		);

	sw_sliders : component nios_ii_base_SW_SLIDERS
		port map (
			clk        => clk_clk,                                                            --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                     --                      reset.reset
			address    => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_readdata,   --                           .readdata
			SW         => sw_sliders_export,                                                  --         external_interface.export
			irq        => irq_mapper_receiver0_irq                                            --                  interrupt.irq
		);

	vga_char_buffer : component nios_ii_base_VGA_Char_Buffer
		port map (
			clk                  => clk_clk,                                                                  --                       clk.clk
			reset                => rst_controller_001_reset_out_reset,                                       --                     reset.reset
			ctrl_address         => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_address(0),   -- avalon_char_control_slave.address
			ctrl_byteenable      => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_byteenable,   --                          .byteenable
			ctrl_chipselect      => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_chipselect,   --                          .chipselect
			ctrl_read            => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_read,         --                          .read
			ctrl_write           => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_write,        --                          .write
			ctrl_writedata       => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_writedata,    --                          .writedata
			ctrl_readdata        => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_readdata,     --                          .readdata
			buf_byteenable       => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_byteenable(0), --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_chipselect,    --                          .chipselect
			buf_read             => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_read,          --                          .read
			buf_write            => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_write,         --                          .write
			buf_writedata        => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_writedata,     --                          .writedata
			buf_readdata         => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_readdata,      --                          .readdata
			buf_waitrequest      => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_waitrequest,   --                          .waitrequest
			buf_address          => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_address,       --                          .address
			stream_ready         => vga_char_buffer_avalon_char_source_ready,                                 --        avalon_char_source.ready
			stream_startofpacket => vga_char_buffer_avalon_char_source_startofpacket,                         --                          .startofpacket
			stream_endofpacket   => vga_char_buffer_avalon_char_source_endofpacket,                           --                          .endofpacket
			stream_valid         => vga_char_buffer_avalon_char_source_valid,                                 --                          .valid
			stream_data          => vga_char_buffer_avalon_char_source_data                                   --                          .data
		);

	vga_controller : component nios_ii_base_VGA_Controller
		port map (
			clk           => vga_pll_vga_clk_clk,                                       --                clk.clk
			reset         => rst_controller_002_reset_out_reset,                        --              reset.reset
			data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                   -- external_interface.export
			VGA_HS        => vga_HS,                                                    --                   .export
			VGA_VS        => vga_VS,                                                    --                   .export
			VGA_BLANK     => vga_BLANK,                                                 --                   .export
			VGA_SYNC      => vga_SYNC,                                                  --                   .export
			VGA_R         => vga_R,                                                     --                   .export
			VGA_G         => vga_G,                                                     --                   .export
			VGA_B         => vga_B                                                      --                   .export
		);

	vga_dual_clock_fifo : component nios_ii_base_VGA_Dual_Clock_FIFO
		port map (
			clk_stream_in            => clk_clk,                                                   --         clock_stream_in.clk
			reset_stream_in          => rst_controller_001_reset_out_reset,                        --         reset_stream_in.reset
			clk_stream_out           => vga_pll_vga_clk_clk,                                       --        clock_stream_out.clk
			reset_stream_out         => rst_controller_002_reset_out_reset,                        --        reset_stream_out.reset
			stream_in_ready          => vga_char_buffer_avalon_char_source_ready,                  --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => vga_char_buffer_avalon_char_source_startofpacket,          --                        .startofpacket
			stream_in_endofpacket    => vga_char_buffer_avalon_char_source_endofpacket,            --                        .endofpacket
			stream_in_valid          => vga_char_buffer_avalon_char_source_valid,                  --                        .valid
			stream_in_data           => vga_char_buffer_avalon_char_source_data,                   --                        .data
			stream_out_ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	vga_pll : component nios_ii_base_VGA_PLL
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => vga_pll_vga_clk_clk,                --      vga_clk.clk
			reset_source_reset => vga_pll_reset_source_reset          -- reset_source.reset
		);

	timer_0 : component nios_ii_base_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	timer_1 : component nios_ii_base_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                      --   irq.irq
		);

	mm_interconnect_0 : component nios_ii_base_mm_interconnect_0
		port map (
			clk_0_clk_clk                                        => clk_clk,                                                                --                                     clk_0_clk.clk
			NIOS_II_Processor_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                         -- NIOS_II_Processor_reset_reset_bridge_in_reset.reset
			VGA_Char_Buffer_reset_reset_bridge_in_reset_reset    => rst_controller_001_reset_out_reset,                                     --   VGA_Char_Buffer_reset_reset_bridge_in_reset.reset
			NIOS_II_Processor_data_master_address                => nios_ii_processor_data_master_address,                                  --                 NIOS_II_Processor_data_master.address
			NIOS_II_Processor_data_master_waitrequest            => nios_ii_processor_data_master_waitrequest,                              --                                              .waitrequest
			NIOS_II_Processor_data_master_byteenable             => nios_ii_processor_data_master_byteenable,                               --                                              .byteenable
			NIOS_II_Processor_data_master_read                   => nios_ii_processor_data_master_read,                                     --                                              .read
			NIOS_II_Processor_data_master_readdata               => nios_ii_processor_data_master_readdata,                                 --                                              .readdata
			NIOS_II_Processor_data_master_write                  => nios_ii_processor_data_master_write,                                    --                                              .write
			NIOS_II_Processor_data_master_writedata              => nios_ii_processor_data_master_writedata,                                --                                              .writedata
			NIOS_II_Processor_data_master_debugaccess            => nios_ii_processor_data_master_debugaccess,                              --                                              .debugaccess
			NIOS_II_Processor_instruction_master_address         => nios_ii_processor_instruction_master_address,                           --          NIOS_II_Processor_instruction_master.address
			NIOS_II_Processor_instruction_master_waitrequest     => nios_ii_processor_instruction_master_waitrequest,                       --                                              .waitrequest
			NIOS_II_Processor_instruction_master_read            => nios_ii_processor_instruction_master_read,                              --                                              .read
			NIOS_II_Processor_instruction_master_readdata        => nios_ii_processor_instruction_master_readdata,                          --                                              .readdata
			HEX_3_avalon_parallel_port_slave_address             => mm_interconnect_0_hex_3_avalon_parallel_port_slave_address,             --              HEX_3_avalon_parallel_port_slave.address
			HEX_3_avalon_parallel_port_slave_write               => mm_interconnect_0_hex_3_avalon_parallel_port_slave_write,               --                                              .write
			HEX_3_avalon_parallel_port_slave_read                => mm_interconnect_0_hex_3_avalon_parallel_port_slave_read,                --                                              .read
			HEX_3_avalon_parallel_port_slave_readdata            => mm_interconnect_0_hex_3_avalon_parallel_port_slave_readdata,            --                                              .readdata
			HEX_3_avalon_parallel_port_slave_writedata           => mm_interconnect_0_hex_3_avalon_parallel_port_slave_writedata,           --                                              .writedata
			HEX_3_avalon_parallel_port_slave_byteenable          => mm_interconnect_0_hex_3_avalon_parallel_port_slave_byteenable,          --                                              .byteenable
			HEX_3_avalon_parallel_port_slave_chipselect          => mm_interconnect_0_hex_3_avalon_parallel_port_slave_chipselect,          --                                              .chipselect
			HEX_7_avalon_parallel_port_slave_address             => mm_interconnect_0_hex_7_avalon_parallel_port_slave_address,             --              HEX_7_avalon_parallel_port_slave.address
			HEX_7_avalon_parallel_port_slave_write               => mm_interconnect_0_hex_7_avalon_parallel_port_slave_write,               --                                              .write
			HEX_7_avalon_parallel_port_slave_read                => mm_interconnect_0_hex_7_avalon_parallel_port_slave_read,                --                                              .read
			HEX_7_avalon_parallel_port_slave_readdata            => mm_interconnect_0_hex_7_avalon_parallel_port_slave_readdata,            --                                              .readdata
			HEX_7_avalon_parallel_port_slave_writedata           => mm_interconnect_0_hex_7_avalon_parallel_port_slave_writedata,           --                                              .writedata
			HEX_7_avalon_parallel_port_slave_byteenable          => mm_interconnect_0_hex_7_avalon_parallel_port_slave_byteenable,          --                                              .byteenable
			HEX_7_avalon_parallel_port_slave_chipselect          => mm_interconnect_0_hex_7_avalon_parallel_port_slave_chipselect,          --                                              .chipselect
			JTAG_UART_avalon_jtag_slave_address                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                  --                   JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                    --                                              .write
			JTAG_UART_avalon_jtag_slave_read                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                     --                                              .read
			JTAG_UART_avalon_jtag_slave_readdata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                 --                                              .readdata
			JTAG_UART_avalon_jtag_slave_writedata                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                --                                              .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,              --                                              .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,               --                                              .chipselect
			LCD_avalon_lcd_slave_address                         => mm_interconnect_0_lcd_avalon_lcd_slave_address,                         --                          LCD_avalon_lcd_slave.address
			LCD_avalon_lcd_slave_write                           => mm_interconnect_0_lcd_avalon_lcd_slave_write,                           --                                              .write
			LCD_avalon_lcd_slave_read                            => mm_interconnect_0_lcd_avalon_lcd_slave_read,                            --                                              .read
			LCD_avalon_lcd_slave_readdata                        => mm_interconnect_0_lcd_avalon_lcd_slave_readdata,                        --                                              .readdata
			LCD_avalon_lcd_slave_writedata                       => mm_interconnect_0_lcd_avalon_lcd_slave_writedata,                       --                                              .writedata
			LCD_avalon_lcd_slave_waitrequest                     => mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest,                     --                                              .waitrequest
			LCD_avalon_lcd_slave_chipselect                      => mm_interconnect_0_lcd_avalon_lcd_slave_chipselect,                      --                                              .chipselect
			LEDS_GREEN_avalon_parallel_port_slave_address        => mm_interconnect_0_leds_green_avalon_parallel_port_slave_address,        --         LEDS_GREEN_avalon_parallel_port_slave.address
			LEDS_GREEN_avalon_parallel_port_slave_write          => mm_interconnect_0_leds_green_avalon_parallel_port_slave_write,          --                                              .write
			LEDS_GREEN_avalon_parallel_port_slave_read           => mm_interconnect_0_leds_green_avalon_parallel_port_slave_read,           --                                              .read
			LEDS_GREEN_avalon_parallel_port_slave_readdata       => mm_interconnect_0_leds_green_avalon_parallel_port_slave_readdata,       --                                              .readdata
			LEDS_GREEN_avalon_parallel_port_slave_writedata      => mm_interconnect_0_leds_green_avalon_parallel_port_slave_writedata,      --                                              .writedata
			LEDS_GREEN_avalon_parallel_port_slave_byteenable     => mm_interconnect_0_leds_green_avalon_parallel_port_slave_byteenable,     --                                              .byteenable
			LEDS_GREEN_avalon_parallel_port_slave_chipselect     => mm_interconnect_0_leds_green_avalon_parallel_port_slave_chipselect,     --                                              .chipselect
			LEDS_RED_avalon_parallel_port_slave_address          => mm_interconnect_0_leds_red_avalon_parallel_port_slave_address,          --           LEDS_RED_avalon_parallel_port_slave.address
			LEDS_RED_avalon_parallel_port_slave_write            => mm_interconnect_0_leds_red_avalon_parallel_port_slave_write,            --                                              .write
			LEDS_RED_avalon_parallel_port_slave_read             => mm_interconnect_0_leds_red_avalon_parallel_port_slave_read,             --                                              .read
			LEDS_RED_avalon_parallel_port_slave_readdata         => mm_interconnect_0_leds_red_avalon_parallel_port_slave_readdata,         --                                              .readdata
			LEDS_RED_avalon_parallel_port_slave_writedata        => mm_interconnect_0_leds_red_avalon_parallel_port_slave_writedata,        --                                              .writedata
			LEDS_RED_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_leds_red_avalon_parallel_port_slave_byteenable,       --                                              .byteenable
			LEDS_RED_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_leds_red_avalon_parallel_port_slave_chipselect,       --                                              .chipselect
			NIOS_II_Processor_debug_mem_slave_address            => mm_interconnect_0_nios_ii_processor_debug_mem_slave_address,            --             NIOS_II_Processor_debug_mem_slave.address
			NIOS_II_Processor_debug_mem_slave_write              => mm_interconnect_0_nios_ii_processor_debug_mem_slave_write,              --                                              .write
			NIOS_II_Processor_debug_mem_slave_read               => mm_interconnect_0_nios_ii_processor_debug_mem_slave_read,               --                                              .read
			NIOS_II_Processor_debug_mem_slave_readdata           => mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata,           --                                              .readdata
			NIOS_II_Processor_debug_mem_slave_writedata          => mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata,          --                                              .writedata
			NIOS_II_Processor_debug_mem_slave_byteenable         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable,         --                                              .byteenable
			NIOS_II_Processor_debug_mem_slave_waitrequest        => mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest,        --                                              .waitrequest
			NIOS_II_Processor_debug_mem_slave_debugaccess        => mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess,        --                                              .debugaccess
			OnChip_Memory_s1_address                             => mm_interconnect_0_onchip_memory_s1_address,                             --                              OnChip_Memory_s1.address
			OnChip_Memory_s1_write                               => mm_interconnect_0_onchip_memory_s1_write,                               --                                              .write
			OnChip_Memory_s1_readdata                            => mm_interconnect_0_onchip_memory_s1_readdata,                            --                                              .readdata
			OnChip_Memory_s1_writedata                           => mm_interconnect_0_onchip_memory_s1_writedata,                           --                                              .writedata
			OnChip_Memory_s1_byteenable                          => mm_interconnect_0_onchip_memory_s1_byteenable,                          --                                              .byteenable
			OnChip_Memory_s1_chipselect                          => mm_interconnect_0_onchip_memory_s1_chipselect,                          --                                              .chipselect
			OnChip_Memory_s1_clken                               => mm_interconnect_0_onchip_memory_s1_clken,                               --                                              .clken
			Pushbuttons_avalon_parallel_port_slave_address       => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address,       --        Pushbuttons_avalon_parallel_port_slave.address
			Pushbuttons_avalon_parallel_port_slave_write         => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write,         --                                              .write
			Pushbuttons_avalon_parallel_port_slave_read          => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read,          --                                              .read
			Pushbuttons_avalon_parallel_port_slave_readdata      => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata,      --                                              .readdata
			Pushbuttons_avalon_parallel_port_slave_writedata     => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata,     --                                              .writedata
			Pushbuttons_avalon_parallel_port_slave_byteenable    => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable,    --                                              .byteenable
			Pushbuttons_avalon_parallel_port_slave_chipselect    => mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect,    --                                              .chipselect
			SW_SLIDERS_avalon_parallel_port_slave_address        => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_address,        --         SW_SLIDERS_avalon_parallel_port_slave.address
			SW_SLIDERS_avalon_parallel_port_slave_write          => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_write,          --                                              .write
			SW_SLIDERS_avalon_parallel_port_slave_read           => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_read,           --                                              .read
			SW_SLIDERS_avalon_parallel_port_slave_readdata       => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_readdata,       --                                              .readdata
			SW_SLIDERS_avalon_parallel_port_slave_writedata      => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_writedata,      --                                              .writedata
			SW_SLIDERS_avalon_parallel_port_slave_byteenable     => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_byteenable,     --                                              .byteenable
			SW_SLIDERS_avalon_parallel_port_slave_chipselect     => mm_interconnect_0_sw_sliders_avalon_parallel_port_slave_chipselect,     --                                              .chipselect
			timer_0_s1_address                                   => mm_interconnect_0_timer_0_s1_address,                                   --                                    timer_0_s1.address
			timer_0_s1_write                                     => mm_interconnect_0_timer_0_s1_write,                                     --                                              .write
			timer_0_s1_readdata                                  => mm_interconnect_0_timer_0_s1_readdata,                                  --                                              .readdata
			timer_0_s1_writedata                                 => mm_interconnect_0_timer_0_s1_writedata,                                 --                                              .writedata
			timer_0_s1_chipselect                                => mm_interconnect_0_timer_0_s1_chipselect,                                --                                              .chipselect
			timer_1_s1_address                                   => mm_interconnect_0_timer_1_s1_address,                                   --                                    timer_1_s1.address
			timer_1_s1_write                                     => mm_interconnect_0_timer_1_s1_write,                                     --                                              .write
			timer_1_s1_readdata                                  => mm_interconnect_0_timer_1_s1_readdata,                                  --                                              .readdata
			timer_1_s1_writedata                                 => mm_interconnect_0_timer_1_s1_writedata,                                 --                                              .writedata
			timer_1_s1_chipselect                                => mm_interconnect_0_timer_1_s1_chipselect,                                --                                              .chipselect
			VGA_Char_Buffer_avalon_char_buffer_slave_address     => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_address,     --      VGA_Char_Buffer_avalon_char_buffer_slave.address
			VGA_Char_Buffer_avalon_char_buffer_slave_write       => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_write,       --                                              .write
			VGA_Char_Buffer_avalon_char_buffer_slave_read        => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_read,        --                                              .read
			VGA_Char_Buffer_avalon_char_buffer_slave_readdata    => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_readdata,    --                                              .readdata
			VGA_Char_Buffer_avalon_char_buffer_slave_writedata   => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_writedata,   --                                              .writedata
			VGA_Char_Buffer_avalon_char_buffer_slave_byteenable  => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_byteenable,  --                                              .byteenable
			VGA_Char_Buffer_avalon_char_buffer_slave_waitrequest => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_waitrequest, --                                              .waitrequest
			VGA_Char_Buffer_avalon_char_buffer_slave_chipselect  => mm_interconnect_0_vga_char_buffer_avalon_char_buffer_slave_chipselect,  --                                              .chipselect
			VGA_Char_Buffer_avalon_char_control_slave_address    => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_address,    --     VGA_Char_Buffer_avalon_char_control_slave.address
			VGA_Char_Buffer_avalon_char_control_slave_write      => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_write,      --                                              .write
			VGA_Char_Buffer_avalon_char_control_slave_read       => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_read,       --                                              .read
			VGA_Char_Buffer_avalon_char_control_slave_readdata   => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_readdata,   --                                              .readdata
			VGA_Char_Buffer_avalon_char_control_slave_writedata  => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_writedata,  --                                              .writedata
			VGA_Char_Buffer_avalon_char_control_slave_byteenable => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_byteenable, --                                              .byteenable
			VGA_Char_Buffer_avalon_char_control_slave_chipselect => mm_interconnect_0_vga_char_buffer_avalon_char_control_slave_chipselect  --                                              .chipselect
		);

	irq_mapper : component nios_ii_base_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			sender_irq    => nios_ii_processor_irq_irq       --    sender.irq
		);

	rst_controller : component nios_ii_base_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                     -- reset_in0.reset
			reset_in1      => nios_ii_processor_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset,              -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,          --          .reset_req
			reset_req_in0  => '0',                                         -- (terminated)
			reset_req_in1  => '0',                                         -- (terminated)
			reset_in2      => '0',                                         -- (terminated)
			reset_req_in2  => '0',                                         -- (terminated)
			reset_in3      => '0',                                         -- (terminated)
			reset_req_in3  => '0',                                         -- (terminated)
			reset_in4      => '0',                                         -- (terminated)
			reset_req_in4  => '0',                                         -- (terminated)
			reset_in5      => '0',                                         -- (terminated)
			reset_req_in5  => '0',                                         -- (terminated)
			reset_in6      => '0',                                         -- (terminated)
			reset_req_in6  => '0',                                         -- (terminated)
			reset_in7      => '0',                                         -- (terminated)
			reset_req_in7  => '0',                                         -- (terminated)
			reset_in8      => '0',                                         -- (terminated)
			reset_req_in8  => '0',                                         -- (terminated)
			reset_in9      => '0',                                         -- (terminated)
			reset_req_in9  => '0',                                         -- (terminated)
			reset_in10     => '0',                                         -- (terminated)
			reset_req_in10 => '0',                                         -- (terminated)
			reset_in11     => '0',                                         -- (terminated)
			reset_req_in11 => '0',                                         -- (terminated)
			reset_in12     => '0',                                         -- (terminated)
			reset_req_in12 => '0',                                         -- (terminated)
			reset_in13     => '0',                                         -- (terminated)
			reset_req_in13 => '0',                                         -- (terminated)
			reset_in14     => '0',                                         -- (terminated)
			reset_req_in14 => '0',                                         -- (terminated)
			reset_in15     => '0',                                         -- (terminated)
			reset_req_in15 => '0'                                          -- (terminated)
		);

	rst_controller_001 : component nios_ii_base_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios_ii_base_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => vga_pll_reset_source_reset,         -- reset_in0.reset
			clk            => vga_pll_vga_clk_clk,                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_ii_base
